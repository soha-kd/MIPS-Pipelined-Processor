library verilog;
use verilog.vl_types.all;
entity MIPS_PP_tb is
end MIPS_PP_tb;
